* test

.include BSS84.mod

.model nmos nmos(level=14, version=4.6.5)
.model pmos pmos(level=14, version=4.6.5)
* dgsb
.model npn npn(level=1)
.model pnp pnp(level=1)
* cbe

V2 vtemp 0 dc 27v
V1 vcc 0 dc 3.3V

X0 0 ctrl sda vtemp BSS84
*M0 0 ctrl sda 0 pmos
*Cload sda 0 0.1u
R34 ctrl vcc 4.7k
R26 sda vcc 1k

V0 ctrl 0 dc 0V pulse(0 3.3V 1m 10u 10u 1m 2m)
