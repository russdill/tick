* test

.include NDC7002N.mod
.include Si7997DP.mod

.model nmos nmos(level=14, version=4.6.5)
.model pmos pmos(level=14, version=4.6.5)
* Drain gate source substrate
* arrow goes to/from source
* dgsb
.model npn npn(level=1)
.model pnp pnp(level=1)
* cbe

V1 vcc 0 dc 5V


R21 ctrl 0 4.7k
X3 n1 ctrl 0 NDC7002N
R20 vcc n1 4.7k
X2a n2 n1 vcc Si7997DP
R19 n2 0 10k
X2b vout n2 vcc Si7997DP
Rload vout 0 100
C30 vout n2 0.1u

V0 ctrl 0 dc 0V pulse(0 3.3V 50m 5m 5m 50m 100m)
